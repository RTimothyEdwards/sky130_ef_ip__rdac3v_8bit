magic
tech sky130A
magscale 1 2
timestamp 1718228761
<< dnwell >>
rect 5855 109 25830 15769
<< nwell >>
rect 5746 15563 25939 15878
rect 5746 315 6061 15563
rect 25624 315 25939 15563
rect 5746 0 25939 315
<< mvnsubdiff >>
rect 5812 15792 25873 15812
rect 5812 15758 5892 15792
rect 25793 15758 25873 15792
rect 5812 15738 25873 15758
rect 5812 15732 5886 15738
rect 5812 146 5832 15732
rect 5866 146 5886 15732
rect 5812 140 5886 146
rect 25799 15732 25873 15738
rect 25799 146 25819 15732
rect 25853 146 25873 15732
rect 25799 140 25873 146
rect 5812 120 25873 140
rect 5812 86 5892 120
rect 25793 86 25873 120
rect 5812 66 25873 86
<< mvnsubdiffcont >>
rect 5892 15758 25793 15792
rect 5832 146 5866 15732
rect 25819 146 25853 15732
rect 5892 86 25793 120
<< locali >>
rect 11990 16746 12216 16820
rect 5832 15758 5892 15792
rect 25793 15758 25853 15792
rect 5832 15732 5866 15758
rect 5832 120 5866 146
rect 25819 15732 25853 15758
rect 25819 120 25853 146
rect 5832 86 5892 120
rect 25793 86 25853 120
<< viali >>
rect 5903 15758 25782 15792
rect 5832 158 5866 15720
rect 25819 156 25853 15720
rect 5903 86 25781 120
<< metal1 >>
rect 1593 16944 12534 17118
rect 1593 15070 1767 16944
rect 4435 16747 4445 16817
rect 4727 16797 4737 16817
rect 11990 16810 12216 16820
rect 11990 16797 11998 16810
rect 4727 16761 11998 16797
rect 4727 16747 4737 16761
rect 11990 16754 11998 16761
rect 12206 16754 12216 16810
rect 11990 16746 12216 16754
rect 5812 15792 25873 15812
rect 5812 15758 5903 15792
rect 25782 15758 25873 15792
rect 5812 15738 25873 15758
rect 5812 15720 5886 15738
rect 1593 15048 1812 15070
rect 1593 14460 1614 15048
rect 1792 14460 1812 15048
rect 1593 14441 1812 14460
rect 4293 13575 4303 13585
rect -200 13539 4303 13575
rect 4293 13523 4303 13539
rect 4523 13523 4533 13585
rect 4545 13135 4597 13136
rect 4440 12927 4545 13135
rect 4597 12927 4610 13135
rect -200 12091 124 12149
rect 4440 11983 4621 12191
rect 4673 11983 4688 12191
rect 4697 11507 4749 11508
rect 4440 11299 4697 11507
rect 4749 11299 4761 11507
rect -200 10463 124 10521
rect 4440 10355 4773 10563
rect 4825 10355 4835 10563
rect 4925 9879 4977 9880
rect 4440 9671 4925 9879
rect 4977 9671 4986 9879
rect -200 8835 124 8893
rect 4440 8727 4849 8935
rect 4901 8727 4913 8935
rect 4440 8051 5057 8251
rect 4440 8043 5077 8051
rect 4770 7843 5077 8043
rect 5129 7843 5142 8051
rect -200 7207 124 7265
rect 4440 7099 5001 7307
rect 5053 7099 5061 7307
rect 5229 6623 5281 6624
rect 4440 6415 5229 6623
rect 5281 6415 5291 6623
rect -200 5579 124 5637
rect 4440 5471 5153 5679
rect 5205 5471 5218 5679
rect 5381 4995 5433 4996
rect 4440 4787 5381 4995
rect 5433 4787 5445 4995
rect -200 3951 124 4009
rect 4440 3843 5305 4051
rect 5357 3843 5370 4051
rect 5533 3487 5585 3488
rect 5108 3367 5533 3487
rect 4440 3280 5533 3367
rect 5585 3280 5597 3487
rect 4440 3160 5335 3280
rect -200 2323 124 2381
rect 4440 2215 5457 2423
rect 5509 2215 5524 2423
rect 5609 1738 5661 1739
rect 4446 1531 5609 1738
rect 5661 1531 5669 1738
rect -200 695 124 753
rect 4440 587 5687 795
rect 5739 587 5747 795
rect 5812 158 5832 15720
rect 5866 158 5886 15720
rect 25799 15720 25873 15738
rect 5957 15628 6185 15659
rect 25799 15651 25819 15720
rect 5957 262 5997 15628
rect 6143 262 6185 15628
rect 25504 15603 25819 15651
rect 7254 1530 7369 1930
rect 24310 1530 24425 1930
rect 6304 841 6354 1459
rect 7204 1443 7210 1530
rect 7413 1443 7419 1530
rect 24260 1443 24266 1530
rect 24469 1443 24475 1530
rect 25325 837 25375 1461
rect 5957 217 6185 262
rect 25504 237 25544 15603
rect 25690 237 25819 15603
rect 25504 209 25819 237
rect 25728 205 25819 209
rect 5812 140 5886 158
rect 25799 156 25819 205
rect 25853 156 25873 15720
rect 25799 140 25873 156
rect 5812 120 25873 140
rect 5812 86 5903 120
rect 25781 86 25873 120
rect 5812 66 25873 86
<< via1 >>
rect 4445 16747 4727 16817
rect 11998 16754 12206 16810
rect 1614 14460 1792 15048
rect 4303 13523 4523 13585
rect 4545 12927 4597 13135
rect 4621 11983 4673 12191
rect 4697 11299 4749 11507
rect 4773 10355 4825 10563
rect 4925 9671 4977 9879
rect 4849 8727 4901 8935
rect 5077 7843 5129 8051
rect 5001 7099 5053 7307
rect 5229 6415 5281 6623
rect 5153 5471 5205 5679
rect 5381 4787 5433 4995
rect 5305 3843 5357 4051
rect 5533 3280 5585 3487
rect 5457 2215 5509 2423
rect 5609 1531 5661 1738
rect 5687 587 5739 795
rect 5997 262 6143 15628
rect 7210 1443 7413 1530
rect 24266 1443 24469 1530
rect 25544 237 25690 15603
<< metal2 >>
rect 16818 21016 17073 21270
rect 15476 17312 15647 17322
rect 12171 17154 13878 17200
rect 15476 17160 15488 17312
rect 15636 17160 15647 17312
rect 4445 16817 4727 16827
rect 12171 16820 12217 17154
rect 14232 17115 14752 17156
rect 15476 17149 15647 17160
rect 4445 16737 4727 16747
rect 11990 16810 12217 16820
rect 11990 16754 11998 16810
rect 12206 16754 12217 16810
rect 11990 16751 12217 16754
rect 12407 16959 14923 17115
rect 12407 16900 12769 16959
rect 13296 16900 13677 16959
rect 14205 16900 14716 16959
rect 14850 16900 14923 16959
rect 12407 16877 14923 16900
rect 11990 16746 12216 16751
rect -200 15048 1811 15070
rect -200 14691 1614 15048
rect -200 14246 597 14539
rect 1432 14460 1614 14691
rect 1792 14460 1811 15048
rect 304 13413 597 14246
rect 843 14300 1222 14327
rect 843 13651 855 14300
rect 1210 13651 1222 14300
rect 843 13407 1222 13651
rect 1432 13411 1811 14460
rect 3643 14300 4022 14327
rect 3643 13651 3652 14300
rect 4007 13651 4022 14300
rect 3643 13410 4022 13651
rect 4477 13595 4513 16737
rect 12407 16387 12434 16877
rect 14904 16387 14923 16877
rect 12407 16363 14923 16387
rect 15791 17046 16480 17140
rect 17396 17046 17814 17140
rect 18596 17046 19014 17140
rect 19796 17046 20214 17140
rect 20996 17046 21414 17140
rect 15791 16883 21414 17046
rect 15791 16288 15815 16883
rect 14958 16286 15815 16288
rect 14951 16230 14960 16286
rect 15016 16283 15815 16286
rect 21395 16283 21414 16883
rect 15016 16230 21414 16283
rect 25148 16878 25734 16901
rect 25148 16294 25182 16878
rect 25705 16294 25734 16878
rect 25148 16262 25734 16294
rect 14958 16228 21414 16230
rect 4553 16119 19417 16155
rect 4303 13585 4523 13595
rect 4303 13513 4523 13523
rect 4553 13143 4589 16119
rect 4629 16043 19297 16079
rect 4545 13135 4597 13143
rect 4545 12921 4597 12927
rect 4553 12916 4589 12921
rect 4629 12197 4665 16043
rect 4705 15967 21552 16003
rect 4621 12191 4673 12197
rect 4621 11976 4673 11983
rect 4629 11961 4665 11976
rect 4705 11515 4741 15967
rect 4781 15891 21431 15927
rect 4697 11507 4749 11515
rect 4697 11293 4749 11299
rect 4705 11282 4741 11293
rect 4781 10570 4817 15891
rect 5957 15634 6185 15659
rect 25504 15651 25732 16262
rect 5957 14139 5977 15634
rect 6162 14831 6185 15634
rect 6248 15603 25732 15651
rect 6248 15500 25544 15603
rect 25422 15363 25544 15500
rect 6162 14606 6249 14831
rect 6162 14139 6185 14606
rect 4773 10563 4825 10570
rect 4773 10349 4825 10355
rect 4781 10340 4817 10349
rect 4857 8942 4893 13978
rect 4933 9887 4969 13978
rect 4925 9879 4977 9887
rect 4925 9665 4977 9671
rect 4933 9662 4969 9665
rect 4849 8935 4901 8942
rect 4849 8721 4901 8727
rect 4857 8710 4893 8721
rect 5009 7314 5045 13978
rect 5085 8059 5121 13978
rect 5077 8051 5129 8059
rect 5077 7837 5129 7843
rect 5001 7307 5053 7314
rect 5001 7093 5053 7099
rect 5009 2367 5045 7093
rect 5085 2108 5121 7837
rect 5161 5686 5197 13978
rect 5237 6631 5273 13978
rect 5229 6623 5281 6631
rect 5229 6409 5281 6415
rect 5237 6400 5273 6409
rect 5153 5679 5205 5686
rect 5153 5465 5205 5471
rect 5161 5458 5197 5465
rect 5313 4058 5349 13978
rect 5389 5003 5425 13978
rect 5381 4995 5433 5003
rect 5381 4781 5433 4787
rect 5389 4644 5425 4781
rect 5305 4051 5357 4058
rect 5305 3837 5357 3843
rect 5313 3830 5349 3837
rect 5465 2430 5501 13978
rect 5541 3495 5577 13978
rect 5533 3487 5585 3495
rect 5533 3274 5585 3280
rect 5541 3139 5577 3274
rect 5457 2423 5509 2430
rect 5457 2209 5509 2215
rect 5465 2200 5501 2209
rect 5617 1746 5653 13978
rect 5609 1738 5661 1746
rect 5609 1525 5661 1531
rect 5693 887 5729 13978
rect 5693 856 5731 887
rect 5695 802 5731 856
rect 5687 795 5739 802
rect 5687 581 5739 587
rect 5695 572 5731 581
rect 5957 262 5997 14139
rect 6143 13324 6185 14139
rect 25504 14081 25544 15363
rect 25428 13856 25544 14081
rect 15125 13497 15207 13553
rect 23653 13497 23736 13553
rect 6143 13099 6249 13324
rect 6143 11817 6185 13099
rect 25504 12574 25544 13856
rect 25431 12349 25544 12574
rect 6143 11592 6252 11817
rect 6143 10310 6185 11592
rect 25504 11067 25544 12349
rect 25428 10842 25544 11067
rect 6143 10085 6252 10310
rect 6143 8803 6185 10085
rect 25504 9560 25544 10842
rect 25429 9335 25544 9560
rect 6143 8578 6250 8803
rect 6143 7296 6185 8578
rect 25504 8053 25544 9335
rect 25431 7828 25544 8053
rect 6143 7071 6250 7296
rect 6143 5789 6185 7071
rect 25504 6546 25544 7828
rect 25427 6321 25544 6546
rect 6143 5564 6255 5789
rect 6143 4282 6185 5564
rect 25504 5039 25544 6321
rect 25428 4814 25544 5039
rect 6143 4057 6250 4282
rect 6143 2775 6185 4057
rect 25504 3532 25544 4814
rect 25429 3307 25544 3532
rect 6143 2550 6257 2775
rect 6143 1268 6185 2550
rect 25504 2025 25544 3307
rect 25428 1800 25544 2025
rect 24502 1543 24552 1630
rect 24693 1543 24702 1630
rect 24502 1530 24589 1543
rect 6937 1443 6946 1530
rect 7087 1443 7210 1530
rect 7413 1443 7419 1530
rect 24260 1443 24266 1530
rect 24469 1443 24589 1530
rect 6143 1043 6259 1268
rect 6143 262 6185 1043
rect 25504 518 25544 1800
rect 5957 217 6185 262
rect 6248 230 6600 380
rect 25431 380 25544 518
rect 6800 237 25544 380
rect 25690 237 25732 15603
rect 6800 230 25732 237
rect 6248 217 25732 230
rect 25504 209 25732 217
<< via2 >>
rect 15488 17160 15636 17312
rect 855 13651 1210 14300
rect 3652 13651 4007 14300
rect 12434 16387 14904 16877
rect 14960 16230 15016 16286
rect 15815 16283 21395 16883
rect 25182 16294 25705 16878
rect 5977 15628 6162 15634
rect 5977 14139 5997 15628
rect 5997 14139 6143 15628
rect 6143 14139 6162 15628
rect 24552 1543 24693 1630
rect 6946 1443 7087 1530
rect 24846 1050 25031 1261
rect 6600 230 6800 387
<< metal3 >>
rect 15476 17312 15647 17322
rect 15476 17160 15488 17312
rect 15636 17160 15647 17312
rect 15476 17149 15647 17160
rect 5352 16877 14937 16891
rect 5352 16387 12434 16877
rect 14904 16678 14937 16877
rect 14904 16618 15144 16678
rect 14904 16387 14937 16618
rect 5352 16366 14937 16387
rect 5352 16090 6194 16366
rect 14955 16286 15021 16291
rect 14955 16230 14960 16286
rect 15016 16230 15021 16286
rect 14955 16225 15021 16230
rect 5352 15927 5374 16090
rect -200 15699 5374 15927
rect 6170 15699 6194 16090
rect -200 15634 6194 15699
rect -200 15253 5977 15634
rect 3639 14987 4324 15006
rect 3639 14396 3655 14987
rect 4309 14396 4324 14987
rect 3639 14364 4324 14396
rect 3639 14308 4323 14364
rect 826 14300 4323 14308
rect 826 13651 855 14300
rect 1210 13651 3652 14300
rect 4007 13651 4323 14300
rect 5948 14139 5977 15253
rect 6162 14139 6194 15634
rect 8562 15546 8622 16024
rect 8688 15546 8748 15944
rect 10694 15546 10754 16177
rect 10820 15546 10880 16094
rect 12826 15546 12886 15946
rect 12952 15546 13012 16018
rect 14958 15546 15018 16225
rect 15084 15546 15144 16618
rect 5948 14113 6194 14139
rect 8819 14030 8879 14600
rect 10951 14033 11011 14601
rect 9158 13769 9495 13829
rect 5942 13765 5948 13767
rect 4916 13705 5948 13765
rect 5942 13703 5948 13705
rect 6186 13765 6192 13767
rect 6186 13705 6195 13765
rect 6186 13703 6192 13705
rect 826 13640 4323 13651
rect 5942 13636 5948 13638
rect 5595 13576 5948 13636
rect 5942 13574 5948 13576
rect 6186 13636 6192 13638
rect 6186 13576 6195 13636
rect 9158 13594 9218 13769
rect 9620 13678 9682 13697
rect 9493 13618 9682 13678
rect 6186 13574 6192 13576
rect 9493 13534 9559 13618
rect 5942 13507 5948 13509
rect 4911 13447 5948 13507
rect 5942 13445 5948 13447
rect 6186 13507 6192 13509
rect 6186 13447 6195 13507
rect 6186 13445 6192 13447
rect 5942 13378 5948 13380
rect 5671 13318 5948 13378
rect 5942 13316 5948 13318
rect 6186 13378 6192 13380
rect 6186 13318 6195 13378
rect 11262 13326 11322 15391
rect 15520 15372 15580 17149
rect 25148 16900 25734 16901
rect 15791 16883 25734 16900
rect 15791 16283 15815 16883
rect 21395 16878 25734 16883
rect 21395 16848 25182 16878
rect 23389 16315 25182 16848
rect 21395 16294 25182 16315
rect 25705 16294 25734 16878
rect 21395 16283 25734 16294
rect 15791 16262 25734 16283
rect 17090 15564 17150 16021
rect 17216 15564 17276 15943
rect 19222 15564 19282 16099
rect 19348 15564 19408 16171
rect 21354 15564 21414 15945
rect 21480 15564 21540 16017
rect 23486 15564 23546 16262
rect 23612 15706 23622 16056
rect 23744 15706 23754 16056
rect 23612 15568 23672 15706
rect 13083 14032 13143 14601
rect 17347 14032 17407 14601
rect 19479 14033 19539 14601
rect 13422 13769 13763 13829
rect 17686 13769 18027 13829
rect 13422 13509 13482 13769
rect 13884 13678 13946 13703
rect 13757 13618 13946 13678
rect 13757 13455 13823 13618
rect 17686 13509 17746 13769
rect 18148 13678 18210 13703
rect 18021 13618 18210 13678
rect 18021 13455 18087 13618
rect 19790 13335 19850 15400
rect 21611 14032 21671 14601
rect 21950 13769 22291 13829
rect 21950 13509 22010 13769
rect 22412 13678 22474 13703
rect 22285 13618 22474 13678
rect 22285 13455 22351 13618
rect 6186 13316 6192 13318
rect 5942 13111 5948 13113
rect 5593 13051 5948 13111
rect 5942 13049 5948 13051
rect 6186 13111 6192 13113
rect 6186 13051 6195 13111
rect 6186 13049 6192 13051
rect 5942 12982 5948 12984
rect 5440 12922 5948 12982
rect 5942 12920 5948 12922
rect 6186 12982 6192 12984
rect 6186 12922 6195 12982
rect 6186 12920 6192 12922
rect 5942 12853 5948 12855
rect 5670 12793 5948 12853
rect 5942 12791 5948 12793
rect 6186 12853 6192 12855
rect 6186 12793 6195 12853
rect 6186 12791 6192 12793
rect 5942 12724 5948 12726
rect 5521 12664 5948 12724
rect 5942 12662 5948 12664
rect 6186 12724 6192 12726
rect 6186 12664 6195 12724
rect 6186 12662 6192 12664
rect 5942 12258 5948 12260
rect 5444 12198 5948 12258
rect 5942 12196 5948 12198
rect 6186 12258 6192 12260
rect 6186 12198 6195 12258
rect 6186 12196 6192 12198
rect 5942 12129 5948 12131
rect 5667 12069 5948 12129
rect 5942 12067 5948 12069
rect 6186 12129 6192 12131
rect 6186 12069 6195 12129
rect 6186 12067 6192 12069
rect 5942 12000 5948 12002
rect 5518 11940 5948 12000
rect 5942 11938 5948 11940
rect 6186 12000 6192 12002
rect 6186 11940 6195 12000
rect 6186 11938 6192 11940
rect 5942 11871 5948 11873
rect 5595 11811 5948 11871
rect 5942 11809 5948 11811
rect 6186 11871 6192 11873
rect 6186 11811 6195 11871
rect 6186 11809 6192 11811
rect 5942 11604 5948 11606
rect 5671 11544 5948 11604
rect 5942 11542 5948 11544
rect 6186 11604 6192 11606
rect 6186 11544 6195 11604
rect 6186 11542 6192 11544
rect 5942 11475 5948 11477
rect 5294 11415 5948 11475
rect 5942 11413 5948 11415
rect 6186 11475 6192 11477
rect 6186 11415 6195 11475
rect 6186 11413 6192 11415
rect 5942 11346 5948 11348
rect 5597 11286 5948 11346
rect 5942 11284 5948 11286
rect 6186 11346 6192 11348
rect 6186 11286 6195 11346
rect 6186 11284 6192 11286
rect 5942 11217 5948 11219
rect 5367 11157 5948 11217
rect 5942 11155 5948 11157
rect 6186 11217 6192 11219
rect 6186 11157 6195 11217
rect 6186 11155 6192 11157
rect 5942 10751 5948 10753
rect 5287 10691 5948 10751
rect 5942 10689 5948 10691
rect 6186 10751 6192 10753
rect 6186 10691 6195 10751
rect 6186 10689 6192 10691
rect 5942 10622 5948 10624
rect 5594 10562 5948 10622
rect 5942 10560 5948 10562
rect 6186 10622 6192 10624
rect 6186 10562 6195 10622
rect 6186 10560 6192 10562
rect 5942 10493 5948 10495
rect 5369 10433 5948 10493
rect 5942 10431 5948 10433
rect 6186 10493 6192 10495
rect 6186 10433 6195 10493
rect 6186 10431 6192 10433
rect 5942 10364 5948 10366
rect 5670 10304 5948 10364
rect 5942 10302 5948 10304
rect 6186 10364 6192 10366
rect 6186 10304 6195 10364
rect 6186 10302 6192 10304
rect 5942 10097 5948 10099
rect 5594 10037 5948 10097
rect 5942 10035 5948 10037
rect 6186 10097 6192 10099
rect 6186 10037 6195 10097
rect 6186 10035 6192 10037
rect 5942 9968 5948 9970
rect 5517 9908 5948 9968
rect 5942 9906 5948 9908
rect 6186 9968 6192 9970
rect 6186 9908 6195 9968
rect 6186 9906 6192 9908
rect 5942 9839 5948 9841
rect 5670 9779 5948 9839
rect 5942 9777 5948 9779
rect 6186 9839 6192 9841
rect 6186 9779 6195 9839
rect 6186 9777 6192 9779
rect 5942 9710 5948 9712
rect 5446 9650 5948 9710
rect 5942 9648 5948 9650
rect 6186 9710 6192 9712
rect 6186 9650 6195 9710
rect 6186 9648 6192 9650
rect 5942 9244 5948 9246
rect 5517 9184 5948 9244
rect 5942 9182 5948 9184
rect 6186 9244 6192 9246
rect 6186 9184 6195 9244
rect 6186 9182 6192 9184
rect 5942 9115 5948 9117
rect 5670 9055 5948 9115
rect 5942 9053 5948 9055
rect 6186 9115 6192 9117
rect 6186 9055 6195 9115
rect 6186 9053 6192 9055
rect 5942 8986 5948 8988
rect 5443 8926 5948 8986
rect 5942 8924 5948 8926
rect 6186 8986 6192 8988
rect 6186 8926 6195 8986
rect 6186 8924 6192 8926
rect 5942 8857 5948 8859
rect 5594 8797 5948 8857
rect 5942 8795 5948 8797
rect 6186 8857 6192 8859
rect 6186 8797 6195 8857
rect 6186 8795 6192 8797
rect 5942 8590 5948 8592
rect 5668 8530 5948 8590
rect 5942 8528 5948 8530
rect 6186 8590 6192 8592
rect 6186 8530 6195 8590
rect 6186 8528 6192 8530
rect 5942 8461 5948 8463
rect 5212 8401 5948 8461
rect 5942 8399 5948 8401
rect 6186 8461 6192 8463
rect 6186 8401 6195 8461
rect 6186 8399 6192 8401
rect 5942 8332 5948 8334
rect 5594 8272 5948 8332
rect 5942 8270 5948 8272
rect 6186 8332 6192 8334
rect 6186 8272 6195 8332
rect 6186 8270 6192 8272
rect 5942 8203 5948 8205
rect 5142 8143 5948 8203
rect 5942 8141 5948 8143
rect 6186 8203 6192 8205
rect 6186 8143 6195 8203
rect 6186 8141 6192 8143
rect 5942 7737 5948 7739
rect 5213 7677 5948 7737
rect 5942 7675 5948 7677
rect 6186 7737 6192 7739
rect 6186 7677 6195 7737
rect 6186 7675 6192 7677
rect 5942 7608 5948 7610
rect 5594 7548 5948 7608
rect 5942 7546 5948 7548
rect 6186 7608 6192 7610
rect 6186 7548 6195 7608
rect 6186 7546 6192 7548
rect 5942 7479 5948 7481
rect 5139 7419 5948 7479
rect 5942 7417 5948 7419
rect 6186 7479 6192 7481
rect 6186 7419 6195 7479
rect 6186 7417 6192 7419
rect 5942 7350 5948 7352
rect 5665 7290 5948 7350
rect 5942 7288 5948 7290
rect 6186 7350 6192 7352
rect 6186 7290 6195 7350
rect 6186 7288 6192 7290
rect 5942 7083 5948 7085
rect 5593 7023 5948 7083
rect 5942 7021 5948 7023
rect 6186 7083 6192 7085
rect 6186 7023 6195 7083
rect 6186 7021 6192 7023
rect 5942 6954 5948 6956
rect 5441 6894 5948 6954
rect 5942 6892 5948 6894
rect 6186 6954 6192 6956
rect 6186 6894 6195 6954
rect 6186 6892 6192 6894
rect 5942 6825 5948 6827
rect 5671 6765 5948 6825
rect 5942 6763 5948 6765
rect 6186 6825 6192 6827
rect 6186 6765 6195 6825
rect 6186 6763 6192 6765
rect 5942 6696 5948 6698
rect 5517 6636 5948 6696
rect 5942 6634 5948 6636
rect 6186 6696 6192 6698
rect 6186 6636 6195 6696
rect 6186 6634 6192 6636
rect 5942 6230 5948 6232
rect 5444 6170 5948 6230
rect 5942 6168 5948 6170
rect 6186 6230 6192 6232
rect 6186 6170 6195 6230
rect 6186 6168 6192 6170
rect 5942 6101 5948 6103
rect 5671 6041 5948 6101
rect 5942 6039 5948 6041
rect 6186 6101 6192 6103
rect 6186 6041 6195 6101
rect 6186 6039 6192 6041
rect 5942 5972 5948 5974
rect 5516 5912 5948 5972
rect 5942 5910 5948 5912
rect 6186 5972 6192 5974
rect 6186 5912 6195 5972
rect 6186 5910 6192 5912
rect 5942 5843 5948 5845
rect 5591 5783 5948 5843
rect 5942 5781 5948 5783
rect 6186 5843 6192 5845
rect 6186 5783 6195 5843
rect 6186 5781 6192 5783
rect 5942 5576 5948 5578
rect 5671 5516 5948 5576
rect 5942 5514 5948 5516
rect 6186 5576 6192 5578
rect 6186 5516 6195 5576
rect 6186 5514 6192 5516
rect 5942 5447 5948 5449
rect 5370 5387 5948 5447
rect 5942 5385 5948 5387
rect 6186 5447 6192 5449
rect 6186 5387 6195 5447
rect 6186 5385 6192 5387
rect 5942 5318 5948 5320
rect 5594 5258 5948 5318
rect 5942 5256 5948 5258
rect 6186 5318 6192 5320
rect 6186 5258 6195 5318
rect 6186 5256 6192 5258
rect 5942 5189 5948 5191
rect 5293 5129 5948 5189
rect 5942 5127 5948 5129
rect 6186 5189 6192 5191
rect 6186 5129 6195 5189
rect 6186 5127 6192 5129
rect 5942 4723 5948 4725
rect 5367 4663 5948 4723
rect 5942 4661 5948 4663
rect 6186 4723 6192 4725
rect 6186 4663 6195 4723
rect 6186 4661 6192 4663
rect 5942 4594 5948 4596
rect 5595 4534 5948 4594
rect 5942 4532 5948 4534
rect 6186 4594 6192 4596
rect 6186 4534 6195 4594
rect 6186 4532 6192 4534
rect 5942 4465 5948 4467
rect 5292 4405 5948 4465
rect 5942 4403 5948 4405
rect 6186 4465 6192 4467
rect 6186 4405 6195 4465
rect 6186 4403 6192 4405
rect 5942 4336 5948 4338
rect 5668 4276 5948 4336
rect 5942 4274 5948 4276
rect 6186 4336 6192 4338
rect 6186 4276 6195 4336
rect 6186 4274 6192 4276
rect 5942 4069 5948 4071
rect 5595 4009 5948 4069
rect 5942 4007 5948 4009
rect 6186 4069 6192 4071
rect 6186 4009 6195 4069
rect 6186 4007 6192 4009
rect 5942 3940 5948 3942
rect 5525 3880 5948 3940
rect 5942 3878 5948 3880
rect 6186 3940 6192 3942
rect 6186 3880 6195 3940
rect 6186 3878 6192 3880
rect 5942 3811 5948 3813
rect 5671 3751 5948 3811
rect 5942 3749 5948 3751
rect 6186 3811 6192 3813
rect 6186 3751 6195 3811
rect 6186 3749 6192 3751
rect 5942 3682 5948 3684
rect 5443 3622 5948 3682
rect 5942 3620 5948 3622
rect 6186 3682 6192 3684
rect 6186 3622 6195 3682
rect 6186 3620 6192 3622
rect 5942 3216 5948 3218
rect 5524 3156 5948 3216
rect 5942 3154 5948 3156
rect 6186 3216 6192 3218
rect 6186 3156 6195 3216
rect 6186 3154 6192 3156
rect 5942 3087 5948 3089
rect 5674 3027 5948 3087
rect 5942 3025 5948 3027
rect 6186 3087 6192 3089
rect 6186 3027 6195 3087
rect 6186 3025 6192 3027
rect 5942 2958 5948 2960
rect 5439 2898 5948 2958
rect 5942 2896 5948 2898
rect 6186 2958 6192 2960
rect 6186 2898 6195 2958
rect 6186 2896 6192 2898
rect 5942 2829 5948 2831
rect 5597 2769 5948 2829
rect 5942 2767 5948 2769
rect 6186 2829 6192 2831
rect 6186 2769 6195 2829
rect 6186 2767 6192 2769
rect 5942 2562 5948 2564
rect 5665 2502 5948 2562
rect 5942 2500 5948 2502
rect 6186 2562 6192 2564
rect 6186 2502 6195 2562
rect 6186 2500 6192 2502
rect 5942 2433 5948 2435
rect 5066 2373 5948 2433
rect 5942 2371 5948 2373
rect 6186 2433 6192 2435
rect 6186 2373 6195 2433
rect 6186 2371 6192 2373
rect 5942 2304 5948 2306
rect 5598 2244 5948 2304
rect 5942 2242 5948 2244
rect 6186 2304 6192 2306
rect 6186 2244 6195 2304
rect 6186 2242 6192 2244
rect 5942 2175 5948 2177
rect 5068 2115 5948 2175
rect 5942 2113 5948 2115
rect 6186 2175 6192 2177
rect 6186 2115 6195 2175
rect 6186 2113 6192 2115
rect 24547 1630 24768 1635
rect 24547 1543 24552 1630
rect 24693 1543 24768 1630
rect 6896 1530 7133 1535
rect 6896 1443 6946 1530
rect 7087 1443 7133 1530
rect 6587 602 6814 643
rect 5516 592 6814 602
rect 5516 188 5523 592
rect 5855 387 6814 592
rect 5855 230 6600 387
rect 6800 230 6814 387
rect 5855 188 6814 230
rect 5516 182 6814 188
rect 6339 -200 6814 182
rect 6896 -200 7133 1443
rect 24547 -200 24768 1543
rect 24837 1261 25039 1268
rect 24837 1050 24846 1261
rect 25031 1050 25039 1261
rect 24837 456 25039 1050
rect 24837 447 25874 456
rect 24837 75 25543 447
rect 25865 75 25874 447
rect 24837 66 25874 75
rect 24837 -200 25197 66
<< via3 >>
rect 5374 15699 6170 16090
rect 3655 14396 4309 14987
rect 5948 13703 6186 13767
rect 5948 13574 6186 13638
rect 5948 13445 6186 13509
rect 5948 13316 6186 13380
rect 15860 16315 21395 16848
rect 21395 16315 23389 16848
rect 23622 15706 23744 16056
rect 5948 13049 6186 13113
rect 5948 12920 6186 12984
rect 5948 12791 6186 12855
rect 5948 12662 6186 12726
rect 5948 12196 6186 12260
rect 5948 12067 6186 12131
rect 5948 11938 6186 12002
rect 5948 11809 6186 11873
rect 5948 11542 6186 11606
rect 5948 11413 6186 11477
rect 5948 11284 6186 11348
rect 5948 11155 6186 11219
rect 5948 10689 6186 10753
rect 5948 10560 6186 10624
rect 5948 10431 6186 10495
rect 5948 10302 6186 10366
rect 5948 10035 6186 10099
rect 5948 9906 6186 9970
rect 5948 9777 6186 9841
rect 5948 9648 6186 9712
rect 5948 9182 6186 9246
rect 5948 9053 6186 9117
rect 5948 8924 6186 8988
rect 5948 8795 6186 8859
rect 5948 8528 6186 8592
rect 5948 8399 6186 8463
rect 5948 8270 6186 8334
rect 5948 8141 6186 8205
rect 5948 7675 6186 7739
rect 5948 7546 6186 7610
rect 5948 7417 6186 7481
rect 5948 7288 6186 7352
rect 5948 7021 6186 7085
rect 5948 6892 6186 6956
rect 5948 6763 6186 6827
rect 5948 6634 6186 6698
rect 5948 6168 6186 6232
rect 5948 6039 6186 6103
rect 5948 5910 6186 5974
rect 5948 5781 6186 5845
rect 5948 5514 6186 5578
rect 5948 5385 6186 5449
rect 5948 5256 6186 5320
rect 5948 5127 6186 5191
rect 5948 4661 6186 4725
rect 5948 4532 6186 4596
rect 5948 4403 6186 4467
rect 5948 4274 6186 4338
rect 5948 4007 6186 4071
rect 5948 3878 6186 3942
rect 5948 3749 6186 3813
rect 5948 3620 6186 3684
rect 5948 3154 6186 3218
rect 5948 3025 6186 3089
rect 5948 2896 6186 2960
rect 5948 2767 6186 2831
rect 5948 2500 6186 2564
rect 5948 2371 6186 2435
rect 5948 2242 6186 2306
rect 5948 2113 6186 2177
rect 5523 188 5855 592
rect 25543 75 25865 447
<< metal4 >>
rect -200 16848 25872 16900
rect -200 16315 15860 16848
rect 23389 16315 25872 16848
rect -200 16280 25872 16315
rect 3639 15000 4324 16280
rect 5351 16090 25875 16109
rect 5351 15699 5374 16090
rect 6170 16056 25875 16090
rect 6170 15706 23622 16056
rect 23744 15706 25875 16056
rect 6170 15699 25875 15706
rect 5351 15683 25875 15699
rect 11261 15391 19851 15451
rect 3632 14987 5869 15000
rect 3632 14396 3655 14987
rect 4309 14396 5869 14987
rect 8962 14685 13005 14745
rect 17484 14685 21527 14745
rect 3632 14380 5869 14396
rect 5517 592 5869 14380
rect 5947 13767 6187 13768
rect 5947 13765 5948 13767
rect 5941 13705 5948 13765
rect 5947 13703 5948 13705
rect 6186 13765 6187 13767
rect 6186 13705 6255 13765
rect 7290 13706 7385 13762
rect 6186 13703 6187 13705
rect 5947 13702 6187 13703
rect 5947 13638 6187 13639
rect 5947 13636 5948 13638
rect 5941 13576 5948 13636
rect 5947 13574 5948 13576
rect 6186 13636 6187 13638
rect 6186 13576 6255 13636
rect 6186 13574 6187 13576
rect 5947 13573 6187 13574
rect 5947 13509 6187 13510
rect 5947 13507 5948 13509
rect 5941 13447 5948 13507
rect 5947 13445 5948 13447
rect 6186 13507 6187 13509
rect 6186 13447 6255 13507
rect 7291 13449 7386 13505
rect 6186 13445 6187 13447
rect 5947 13444 6187 13445
rect 5947 13380 6187 13381
rect 5947 13378 5948 13380
rect 5941 13318 5948 13378
rect 5947 13316 5948 13318
rect 6186 13378 6187 13380
rect 6186 13318 6255 13378
rect 6186 13316 6187 13318
rect 5947 13315 6187 13316
rect 7741 13192 9733 13252
rect 10785 13192 11172 13252
rect 12001 13192 13993 13252
rect 16268 13192 18260 13252
rect 19313 13192 19700 13252
rect 20535 13192 22527 13252
rect 5947 13113 6187 13114
rect 5947 13111 5948 13113
rect 5941 13051 5948 13111
rect 5947 13049 5948 13051
rect 6186 13111 6187 13113
rect 6186 13051 6255 13111
rect 6186 13049 6187 13051
rect 5947 13048 6187 13049
rect 5947 12984 6187 12985
rect 5947 12982 5948 12984
rect 5941 12922 5948 12982
rect 5947 12920 5948 12922
rect 6186 12982 6187 12984
rect 6186 12922 6255 12982
rect 6186 12920 6187 12922
rect 5947 12919 6187 12920
rect 5947 12855 6187 12856
rect 5947 12853 5948 12855
rect 5941 12793 5948 12853
rect 5947 12791 5948 12793
rect 6186 12853 6187 12855
rect 6186 12793 6255 12853
rect 6186 12791 6187 12793
rect 5947 12790 6187 12791
rect 5947 12726 6187 12727
rect 5947 12724 5948 12726
rect 5941 12664 5948 12724
rect 5947 12662 5948 12664
rect 6186 12724 6187 12726
rect 6186 12664 6255 12724
rect 6186 12662 6187 12664
rect 5947 12661 6187 12662
rect 5947 12260 6187 12261
rect 5947 12258 5948 12260
rect 5941 12198 5948 12258
rect 5947 12196 5948 12198
rect 6186 12258 6187 12260
rect 6186 12198 6255 12258
rect 6186 12196 6187 12198
rect 5947 12195 6187 12196
rect 5947 12131 6187 12132
rect 5947 12129 5948 12131
rect 5941 12069 5948 12129
rect 5947 12067 5948 12069
rect 6186 12129 6187 12131
rect 6186 12069 6255 12129
rect 6186 12067 6187 12069
rect 5947 12066 6187 12067
rect 5947 12002 6187 12003
rect 5947 12000 5948 12002
rect 5941 11940 5948 12000
rect 5947 11938 5948 11940
rect 6186 12000 6187 12002
rect 6186 11940 6255 12000
rect 6186 11938 6187 11940
rect 5947 11937 6187 11938
rect 5947 11873 6187 11874
rect 5947 11871 5948 11873
rect 5941 11811 5948 11871
rect 5947 11809 5948 11811
rect 6186 11871 6187 11873
rect 6186 11811 6255 11871
rect 6186 11809 6187 11811
rect 5947 11808 6187 11809
rect 5947 11606 6187 11607
rect 5947 11604 5948 11606
rect 5941 11544 5948 11604
rect 5947 11542 5948 11544
rect 6186 11604 6187 11606
rect 6186 11544 6255 11604
rect 6186 11542 6187 11544
rect 5947 11541 6187 11542
rect 5947 11477 6187 11478
rect 5947 11475 5948 11477
rect 5941 11415 5948 11475
rect 5947 11413 5948 11415
rect 6186 11475 6187 11477
rect 6186 11415 6255 11475
rect 6186 11413 6187 11415
rect 5947 11412 6187 11413
rect 5947 11348 6187 11349
rect 5947 11346 5948 11348
rect 5941 11286 5948 11346
rect 5947 11284 5948 11286
rect 6186 11346 6187 11348
rect 6186 11286 6255 11346
rect 6186 11284 6187 11286
rect 5947 11283 6187 11284
rect 5947 11219 6187 11220
rect 5947 11217 5948 11219
rect 5941 11157 5948 11217
rect 5947 11155 5948 11157
rect 6186 11217 6187 11219
rect 6186 11157 6255 11217
rect 6186 11155 6187 11157
rect 5947 11154 6187 11155
rect 5947 10753 6187 10754
rect 5947 10751 5948 10753
rect 5941 10691 5948 10751
rect 5947 10689 5948 10691
rect 6186 10751 6187 10753
rect 6186 10691 6255 10751
rect 6186 10689 6187 10691
rect 5947 10688 6187 10689
rect 5947 10624 6187 10625
rect 5947 10622 5948 10624
rect 5941 10562 5948 10622
rect 5947 10560 5948 10562
rect 6186 10622 6187 10624
rect 6186 10562 6255 10622
rect 6186 10560 6187 10562
rect 5947 10559 6187 10560
rect 5947 10495 6187 10496
rect 5947 10493 5948 10495
rect 5941 10433 5948 10493
rect 5947 10431 5948 10433
rect 6186 10493 6187 10495
rect 6186 10433 6255 10493
rect 6186 10431 6187 10433
rect 5947 10430 6187 10431
rect 5947 10366 6187 10367
rect 5947 10364 5948 10366
rect 5941 10304 5948 10364
rect 5947 10302 5948 10304
rect 6186 10364 6187 10366
rect 6186 10304 6255 10364
rect 6186 10302 6187 10304
rect 5947 10301 6187 10302
rect 5947 10099 6187 10100
rect 5947 10097 5948 10099
rect 5941 10037 5948 10097
rect 5947 10035 5948 10037
rect 6186 10097 6187 10099
rect 6186 10037 6255 10097
rect 6186 10035 6187 10037
rect 5947 10034 6187 10035
rect 5947 9970 6187 9971
rect 5947 9968 5948 9970
rect 5941 9908 5948 9968
rect 5947 9906 5948 9908
rect 6186 9968 6187 9970
rect 6186 9908 6255 9968
rect 6186 9906 6187 9908
rect 5947 9905 6187 9906
rect 5947 9841 6187 9842
rect 5947 9839 5948 9841
rect 5941 9779 5948 9839
rect 5947 9777 5948 9779
rect 6186 9839 6187 9841
rect 6186 9779 6255 9839
rect 6186 9777 6187 9779
rect 5947 9776 6187 9777
rect 5947 9712 6187 9713
rect 5947 9710 5948 9712
rect 5941 9650 5948 9710
rect 5947 9648 5948 9650
rect 6186 9710 6187 9712
rect 6186 9650 6255 9710
rect 6186 9648 6187 9650
rect 5947 9647 6187 9648
rect 5947 9246 6187 9247
rect 5947 9244 5948 9246
rect 5941 9184 5948 9244
rect 5947 9182 5948 9184
rect 6186 9244 6187 9246
rect 6186 9184 6255 9244
rect 6186 9182 6187 9184
rect 5947 9181 6187 9182
rect 5947 9117 6187 9118
rect 5947 9115 5948 9117
rect 5941 9055 5948 9115
rect 5947 9053 5948 9055
rect 6186 9115 6187 9117
rect 6186 9055 6255 9115
rect 6186 9053 6187 9055
rect 5947 9052 6187 9053
rect 5947 8988 6187 8989
rect 5947 8986 5948 8988
rect 5941 8926 5948 8986
rect 5947 8924 5948 8926
rect 6186 8986 6187 8988
rect 6186 8926 6255 8986
rect 6186 8924 6187 8926
rect 5947 8923 6187 8924
rect 5947 8859 6187 8860
rect 5947 8857 5948 8859
rect 5941 8797 5948 8857
rect 5947 8795 5948 8797
rect 6186 8857 6187 8859
rect 6186 8797 6255 8857
rect 6186 8795 6187 8797
rect 5947 8794 6187 8795
rect 5947 8592 6187 8593
rect 5947 8590 5948 8592
rect 5941 8530 5948 8590
rect 5947 8528 5948 8530
rect 6186 8590 6187 8592
rect 6186 8530 6255 8590
rect 6186 8528 6187 8530
rect 5947 8527 6187 8528
rect 5947 8463 6187 8464
rect 5947 8461 5948 8463
rect 5941 8401 5948 8461
rect 5947 8399 5948 8401
rect 6186 8461 6187 8463
rect 6186 8401 6255 8461
rect 6186 8399 6187 8401
rect 5947 8398 6187 8399
rect 5947 8334 6187 8335
rect 5947 8332 5948 8334
rect 5941 8272 5948 8332
rect 5947 8270 5948 8272
rect 6186 8332 6187 8334
rect 6186 8272 6255 8332
rect 6186 8270 6187 8272
rect 5947 8269 6187 8270
rect 5947 8205 6187 8206
rect 5947 8203 5948 8205
rect 5941 8143 5948 8203
rect 5947 8141 5948 8143
rect 6186 8203 6187 8205
rect 6186 8143 6255 8203
rect 6186 8141 6187 8143
rect 5947 8140 6187 8141
rect 5947 7739 6187 7740
rect 5947 7737 5948 7739
rect 5941 7677 5948 7737
rect 5947 7675 5948 7677
rect 6186 7737 6187 7739
rect 6186 7677 6255 7737
rect 6186 7675 6187 7677
rect 5947 7674 6187 7675
rect 5947 7610 6187 7611
rect 5947 7608 5948 7610
rect 5941 7548 5948 7608
rect 5947 7546 5948 7548
rect 6186 7608 6187 7610
rect 6186 7548 6255 7608
rect 6186 7546 6187 7548
rect 5947 7545 6187 7546
rect 5947 7481 6187 7482
rect 5947 7479 5948 7481
rect 5941 7419 5948 7479
rect 5947 7417 5948 7419
rect 6186 7479 6187 7481
rect 6186 7419 6255 7479
rect 6186 7417 6187 7419
rect 5947 7416 6187 7417
rect 5947 7352 6187 7353
rect 5947 7350 5948 7352
rect 5941 7290 5948 7350
rect 5947 7288 5948 7290
rect 6186 7350 6187 7352
rect 6186 7290 6255 7350
rect 6186 7288 6187 7290
rect 5947 7287 6187 7288
rect 5947 7085 6187 7086
rect 5947 7083 5948 7085
rect 5941 7023 5948 7083
rect 5947 7021 5948 7023
rect 6186 7083 6187 7085
rect 6186 7023 6255 7083
rect 6186 7021 6187 7023
rect 5947 7020 6187 7021
rect 5947 6956 6187 6957
rect 5947 6954 5948 6956
rect 5941 6894 5948 6954
rect 5947 6892 5948 6894
rect 6186 6954 6187 6956
rect 6186 6894 6255 6954
rect 6186 6892 6187 6894
rect 5947 6891 6187 6892
rect 5947 6827 6187 6828
rect 5947 6825 5948 6827
rect 5941 6765 5948 6825
rect 5947 6763 5948 6765
rect 6186 6825 6187 6827
rect 6186 6765 6255 6825
rect 6186 6763 6187 6765
rect 5947 6762 6187 6763
rect 5947 6698 6187 6699
rect 5947 6696 5948 6698
rect 5941 6636 5948 6696
rect 5947 6634 5948 6636
rect 6186 6696 6187 6698
rect 6186 6636 6255 6696
rect 6186 6634 6187 6636
rect 5947 6633 6187 6634
rect 5947 6232 6187 6233
rect 5947 6230 5948 6232
rect 5941 6170 5948 6230
rect 5947 6168 5948 6170
rect 6186 6230 6187 6232
rect 6186 6170 6255 6230
rect 6186 6168 6187 6170
rect 5947 6167 6187 6168
rect 5947 6103 6187 6104
rect 5947 6101 5948 6103
rect 5941 6041 5948 6101
rect 5947 6039 5948 6041
rect 6186 6101 6187 6103
rect 6186 6041 6255 6101
rect 6186 6039 6187 6041
rect 5947 6038 6187 6039
rect 5947 5974 6187 5975
rect 5947 5972 5948 5974
rect 5941 5912 5948 5972
rect 5947 5910 5948 5912
rect 6186 5972 6187 5974
rect 6186 5912 6255 5972
rect 6186 5910 6187 5912
rect 5947 5909 6187 5910
rect 5947 5845 6187 5846
rect 5947 5843 5948 5845
rect 5941 5783 5948 5843
rect 5947 5781 5948 5783
rect 6186 5843 6187 5845
rect 6186 5783 6255 5843
rect 6186 5781 6187 5783
rect 5947 5780 6187 5781
rect 5947 5578 6187 5579
rect 5947 5576 5948 5578
rect 5941 5516 5948 5576
rect 5947 5514 5948 5516
rect 6186 5576 6187 5578
rect 6186 5516 6255 5576
rect 6186 5514 6187 5516
rect 5947 5513 6187 5514
rect 5947 5449 6187 5450
rect 5947 5447 5948 5449
rect 5941 5387 5948 5447
rect 5947 5385 5948 5387
rect 6186 5447 6187 5449
rect 6186 5387 6255 5447
rect 6186 5385 6187 5387
rect 5947 5384 6187 5385
rect 5947 5320 6187 5321
rect 5947 5318 5948 5320
rect 5941 5258 5948 5318
rect 5947 5256 5948 5258
rect 6186 5318 6187 5320
rect 6186 5258 6255 5318
rect 6186 5256 6187 5258
rect 5947 5255 6187 5256
rect 5947 5191 6187 5192
rect 5947 5189 5948 5191
rect 5941 5129 5948 5189
rect 5947 5127 5948 5129
rect 6186 5189 6187 5191
rect 6186 5129 6255 5189
rect 6186 5127 6187 5129
rect 5947 5126 6187 5127
rect 5947 4725 6187 4726
rect 5947 4723 5948 4725
rect 5941 4663 5948 4723
rect 5947 4661 5948 4663
rect 6186 4723 6187 4725
rect 6186 4663 6255 4723
rect 6186 4661 6187 4663
rect 5947 4660 6187 4661
rect 5947 4596 6187 4597
rect 5947 4594 5948 4596
rect 5941 4534 5948 4594
rect 5947 4532 5948 4534
rect 6186 4594 6187 4596
rect 6186 4534 6255 4594
rect 6186 4532 6187 4534
rect 5947 4531 6187 4532
rect 5947 4467 6187 4468
rect 5947 4465 5948 4467
rect 5941 4405 5948 4465
rect 5947 4403 5948 4405
rect 6186 4465 6187 4467
rect 6186 4405 6255 4465
rect 6186 4403 6187 4405
rect 5947 4402 6187 4403
rect 5947 4338 6187 4339
rect 5947 4336 5948 4338
rect 5941 4276 5948 4336
rect 5947 4274 5948 4276
rect 6186 4336 6187 4338
rect 6186 4276 6255 4336
rect 6186 4274 6187 4276
rect 5947 4273 6187 4274
rect 5947 4071 6187 4072
rect 5947 4069 5948 4071
rect 5941 4009 5948 4069
rect 5947 4007 5948 4009
rect 6186 4069 6187 4071
rect 6186 4009 6255 4069
rect 6186 4007 6187 4009
rect 5947 4006 6187 4007
rect 5947 3942 6187 3943
rect 5947 3940 5948 3942
rect 5941 3880 5948 3940
rect 5947 3878 5948 3880
rect 6186 3940 6187 3942
rect 6186 3880 6255 3940
rect 6186 3878 6187 3880
rect 5947 3877 6187 3878
rect 5947 3813 6187 3814
rect 5947 3811 5948 3813
rect 5941 3751 5948 3811
rect 5947 3749 5948 3751
rect 6186 3811 6187 3813
rect 6186 3751 6255 3811
rect 6186 3749 6187 3751
rect 5947 3748 6187 3749
rect 5947 3684 6187 3685
rect 5947 3682 5948 3684
rect 5941 3622 5948 3682
rect 5947 3620 5948 3622
rect 6186 3682 6187 3684
rect 6186 3622 6255 3682
rect 6186 3620 6187 3622
rect 5947 3619 6187 3620
rect 5947 3218 6187 3219
rect 5947 3216 5948 3218
rect 5941 3156 5948 3216
rect 5947 3154 5948 3156
rect 6186 3216 6187 3218
rect 6186 3156 6255 3216
rect 6186 3154 6187 3156
rect 5947 3153 6187 3154
rect 5947 3089 6187 3090
rect 5947 3087 5948 3089
rect 5941 3027 5948 3087
rect 5947 3025 5948 3027
rect 6186 3087 6187 3089
rect 6186 3027 6255 3087
rect 6186 3025 6187 3027
rect 5947 3024 6187 3025
rect 5947 2960 6187 2961
rect 5947 2958 5948 2960
rect 5941 2898 5948 2958
rect 5947 2896 5948 2898
rect 6186 2958 6187 2960
rect 6186 2898 6255 2958
rect 6186 2896 6187 2898
rect 5947 2895 6187 2896
rect 5947 2831 6187 2832
rect 5947 2829 5948 2831
rect 5941 2769 5948 2829
rect 5947 2767 5948 2769
rect 6186 2829 6187 2831
rect 6186 2769 6255 2829
rect 6186 2767 6187 2769
rect 5947 2766 6187 2767
rect 5947 2564 6187 2565
rect 5947 2562 5948 2564
rect 5941 2502 5948 2562
rect 5947 2500 5948 2502
rect 6186 2562 6187 2564
rect 6186 2502 6255 2562
rect 6186 2500 6187 2502
rect 5947 2499 6187 2500
rect 5947 2435 6187 2436
rect 5947 2433 5948 2435
rect 5941 2373 5948 2433
rect 5947 2371 5948 2373
rect 6186 2433 6187 2435
rect 6186 2373 6255 2433
rect 6186 2371 6187 2373
rect 5947 2370 6187 2371
rect 5947 2306 6187 2307
rect 5947 2304 5948 2306
rect 5941 2244 5948 2304
rect 5947 2242 5948 2244
rect 6186 2304 6187 2306
rect 6186 2244 6255 2304
rect 6186 2242 6187 2244
rect 5947 2241 6187 2242
rect 5947 2177 6187 2178
rect 5947 2175 5948 2177
rect 5941 2115 5948 2175
rect 5947 2113 5948 2115
rect 6186 2175 6187 2177
rect 6186 2115 6255 2175
rect 6186 2113 6187 2115
rect 5947 2112 6187 2113
rect 5517 188 5523 592
rect 5855 188 5869 592
rect 5517 66 5869 188
rect 25534 447 25875 15683
rect 25534 75 25543 447
rect 25865 75 25875 447
rect 25534 66 25875 75
use dac_3v_column  dac_3v_column_0
array 0 7 2132 0 0 15271
timestamp 1653060931
transform 1 0 7331 0 1 322
box -20 -7 1049 15264
use dac_3v_column_dummy  dac_3v_column_dummy_0
timestamp 1653061945
transform 1 0 6266 0 1 322
box -18 -7 1049 15272
use dac_3v_column_dummy  dac_3v_column_dummy_1
timestamp 1653061945
transform 1 0 24386 0 1 322
box -18 -7 1049 15272
use dac_3v_column_odd  dac_3v_column_odd_0
array 0 7 2132 0 0 15270
timestamp 1653060931
transform 1 0 8398 0 1 322
box -20 -7 1049 15263
use follower_amp  follower_amp_0 ../dependencies/sky130_ef_ip__samplehold/mag
timestamp 1718228583
transform 0 1 12491 1 0 16882
box 0 0 4377 11129
use level_shifter_array  level_shifter_array_0
timestamp 1652995732
transform 1 0 23 0 1 312
box -23 -10 4908 13105
use m2m3contact  m2m3contact_0
timestamp 1652924542
transform 0 1 4224 -1 0 2458
box 276 844 350 997
use m2m3contact  m2m3contact_1
timestamp 1652924542
transform 0 1 4756 -1 0 2586
box 276 844 350 997
use m2m3contact  m2m3contact_2
timestamp 1652924542
transform 0 1 4831 -1 0 2845
box 276 844 350 997
use m2m3contact  m2m3contact_3
timestamp 1652924542
transform 0 1 4679 -1 0 3499
box 276 844 350 997
use m2m3contact  m2m3contact_4
timestamp 1652924542
transform 0 1 4604 -1 0 3241
box 276 844 350 997
use m2m3contact  m2m3contact_5
timestamp 1652924542
transform 0 1 4832 -1 0 4094
box 276 844 350 997
use m2m3contact  m2m3contact_6
timestamp 1652924542
transform 0 1 4755 -1 0 4353
box 276 844 350 997
use m2m3contact  m2m3contact_7
timestamp 1652924542
transform 0 1 4756 -1 0 5601
box 276 844 350 997
use m2m3contact  m2m3contact_8
timestamp 1652924542
transform 0 1 4831 -1 0 5860
box 276 844 350 997
use m2m3contact  m2m3contact_9
timestamp 1652924542
transform 0 1 4452 -1 0 4748
box 276 844 350 997
use m2m3contact  m2m3contact_10
timestamp 1652924542
transform 0 1 4527 -1 0 5006
box 276 844 350 997
use m2m3contact  m2m3contact_11
timestamp 1652924542
transform 0 1 4756 -1 0 8615
box 276 844 350 997
use m2m3contact  m2m3contact_12
timestamp 1652924542
transform 0 1 4831 -1 0 8874
box 276 844 350 997
use m2m3contact  m2m3contact_13
timestamp 1652924542
transform 0 1 4756 -1 0 11629
box 276 844 350 997
use m2m3contact  m2m3contact_14
timestamp 1652924542
transform 0 1 4831 -1 0 11888
box 276 844 350 997
use m2m3contact  m2m3contact_15
timestamp 1652924542
transform 0 1 4755 -1 0 7367
box 276 844 350 997
use m2m3contact  m2m3contact_16
timestamp 1652924542
transform 0 1 4832 -1 0 7108
box 276 844 350 997
use m2m3contact  m2m3contact_17
timestamp 1652924542
transform 0 1 4755 -1 0 10381
box 276 844 350 997
use m2m3contact  m2m3contact_18
timestamp 1652924542
transform 0 1 4832 -1 0 10122
box 276 844 350 997
use m2m3contact  m2m3contact_19
timestamp 1652924542
transform 0 1 4755 -1 0 13395
box 276 844 350 997
use m2m3contact  m2m3contact_20
timestamp 1652924542
transform 0 1 4832 -1 0 13136
box 276 844 350 997
use m2m3contact  m2m3contact_21
timestamp 1652924542
transform 0 1 4680 -1 0 6255
box 276 844 350 997
use m2m3contact  m2m3contact_22
timestamp 1652924542
transform 0 1 4603 -1 0 6513
box 276 844 350 997
use m2m3contact  m2m3contact_23
timestamp 1652924542
transform 0 1 4300 -1 0 7762
box 276 844 350 997
use m2m3contact  m2m3contact_24
timestamp 1652924542
transform 0 1 4375 -1 0 8020
box 276 844 350 997
use m2m3contact  m2m3contact_25
timestamp 1652924542
transform 0 1 4604 -1 0 9269
box 276 844 350 997
use m2m3contact  m2m3contact_26
timestamp 1652924542
transform 0 1 4679 -1 0 9527
box 276 844 350 997
use m2m3contact  m2m3contact_27
timestamp 1652924542
transform 0 1 4528 -1 0 10776
box 276 844 350 997
use m2m3contact  m2m3contact_28
timestamp 1652924542
transform 0 1 4451 -1 0 11034
box 276 844 350 997
use m2m3contact  m2m3contact_29
timestamp 1652924542
transform 0 1 4680 -1 0 12283
box 276 844 350 997
use m2m3contact  m2m3contact_30
timestamp 1652924542
transform 0 1 4603 -1 0 12541
box 276 844 350 997
use m2m3contact  m2m3contact_31
timestamp 1652924542
transform 0 1 3996 -1 0 13790
box 276 844 350 997
use m2m3contact  m2m3contact_32
timestamp 1652924542
transform 0 1 4071 -1 0 14048
box 276 844 350 997
use m2m3contact  m2m3contact_33
timestamp 1652924542
transform 0 1 4148 -1 0 2716
box 276 844 350 997
use m2m3contact  m2m3contact_34
timestamp 1652924542
transform 0 1 4756 -1 0 3112
box 276 844 350 997
use m2m3contact  m2m3contact_35
timestamp 1652924542
transform 0 1 4832 -1 0 3370
box 276 844 350 997
use m2m3contact  m2m3contact_36
timestamp 1652924542
transform 0 1 4832 -1 0 4619
box 276 844 350 997
use m2m3contact  m2m3contact_37
timestamp 1652924542
transform 0 1 4756 -1 0 4877
box 276 844 350 997
use m2m3contact  m2m3contact_38
timestamp 1652924542
transform 0 1 4832 -1 0 7633
box 276 844 350 997
use m2m3contact  m2m3contact_39
timestamp 1652924542
transform 0 1 4756 -1 0 7891
box 276 844 350 997
use m2m3contact  m2m3contact_40
timestamp 1652924542
transform 0 1 4832 -1 0 10647
box 276 844 350 997
use m2m3contact  m2m3contact_41
timestamp 1652924542
transform 0 1 4756 -1 0 10905
box 276 844 350 997
use m2m3contact  m2m3contact_42
timestamp 1652924542
transform 0 1 4832 -1 0 13661
box 276 844 350 997
use m2m3contact  m2m3contact_43
timestamp 1652924542
transform 0 1 4756 -1 0 13919
box 276 844 350 997
use m2m3contact  m2m3contact_44
timestamp 1652924542
transform 0 1 4756 -1 0 6126
box 276 844 350 997
use m2m3contact  m2m3contact_45
timestamp 1652924542
transform 0 1 4832 -1 0 6384
box 276 844 350 997
use m2m3contact  m2m3contact_46
timestamp 1652924542
transform 0 1 4756 -1 0 9140
box 276 844 350 997
use m2m3contact  m2m3contact_47
timestamp 1652924542
transform 0 1 4832 -1 0 9398
box 276 844 350 997
use m2m3contact  m2m3contact_48
timestamp 1652924542
transform 0 1 4756 -1 0 12154
box 276 844 350 997
use m2m3contact  m2m3contact_49
timestamp 1652924542
transform 0 1 4832 -1 0 12412
box 276 844 350 997
use m2m3contact  m2m3contact_50
timestamp 1652924542
transform 0 1 4604 -1 0 3965
box 276 844 350 997
use m2m3contact  m2m3contact_51
timestamp 1652924542
transform 0 1 4680 -1 0 4223
box 276 844 350 997
use m2m3contact  m2m3contact_52
timestamp 1652924542
transform 0 1 4452 -1 0 5472
box 276 844 350 997
use m2m3contact  m2m3contact_53
timestamp 1652924542
transform 0 1 4528 -1 0 5730
box 276 844 350 997
use m2m3contact  m2m3contact_54
timestamp 1652924542
transform 0 1 4680 -1 0 6979
box 276 844 350 997
use m2m3contact  m2m3contact_55
timestamp 1652924542
transform 0 1 4604 -1 0 7237
box 276 844 350 997
use m2m3contact  m2m3contact_56
timestamp 1652924542
transform 0 1 4300 -1 0 8486
box 276 844 350 997
use m2m3contact  m2m3contact_57
timestamp 1652924542
transform 0 1 4376 -1 0 8744
box 276 844 350 997
use m2m3contact  m2m3contact_58
timestamp 1652924542
transform 0 1 4604 -1 0 9993
box 276 844 350 997
use m2m3contact  m2m3contact_59
timestamp 1652924542
transform 0 1 4680 -1 0 10251
box 276 844 350 997
use m2m3contact  m2m3contact_60
timestamp 1652924542
transform 0 1 4528 -1 0 11500
box 276 844 350 997
use m2m3contact  m2m3contact_61
timestamp 1652924542
transform 0 1 4452 -1 0 11758
box 276 844 350 997
use m2m3contact  m2m3contact_62
timestamp 1652924542
transform 0 1 4604 -1 0 13265
box 276 844 350 997
use m2m3contact  m2m3contact_63
timestamp 1652924542
transform 0 1 4680 -1 0 13007
box 276 844 350 997
use m2m3contact  m2m3contact_64
timestamp 1652924542
transform 1 0 8405 0 1 15028
box 276 844 350 997
use m2m3contact  m2m3contact_65
timestamp 1652924542
transform 1 0 8279 0 1 15106
box 276 844 350 997
use m2m3contact  m2m3contact_66
timestamp 1652924542
transform 1 0 10411 0 1 15258
box 276 844 350 997
use m2m3contact  m2m3contact_67
timestamp 1652924542
transform 1 0 10537 0 1 15180
box 276 844 350 997
use m2m3contact  m2m3contact_68
timestamp 1652924542
transform 1 0 12543 0 1 15030
box 276 844 350 997
use m2m3contact  m2m3contact_69
timestamp 1652924542
transform 1 0 12669 0 1 15104
box 276 844 350 997
use m2m3contact  m2m3contact_72
timestamp 1652924542
transform 1 0 16807 0 1 15106
box 276 844 350 997
use m2m3contact  m2m3contact_73
timestamp 1652924542
transform 1 0 16933 0 1 15028
box 276 844 350 997
use m2m3contact  m2m3contact_74
timestamp 1652924542
transform 1 0 18939 0 1 15182
box 276 844 350 997
use m2m3contact  m2m3contact_75
timestamp 1652924542
transform 1 0 19065 0 -1 17017
box 276 844 350 997
use m2m3contact  m2m3contact_76
timestamp 1652924542
transform 1 0 21071 0 1 15030
box 276 844 350 997
use m2m3contact  m2m3contact_77
timestamp 1652924542
transform 1 0 21197 0 1 15104
box 276 844 350 997
use m3m4contact  m3m4contact_0
timestamp 1652924542
transform -1 0 7257 0 1 6239
box -258 7458 -104 7613
use m3m4contact  m3m4contact_1
timestamp 1652924542
transform -1 0 7257 0 1 5981
box -258 7458 -104 7613
use m3m4contact  m3m4contact_2
timestamp 1652924542
transform -1 0 11521 0 1 6239
box -258 7458 -104 7613
use m3m4contact  m3m4contact_3
timestamp 1652924542
transform -1 0 11521 0 1 5981
box -258 7458 -104 7613
use m3m4contact  m3m4contact_4
timestamp 1652924542
transform -1 0 15785 0 1 6239
box -258 7458 -104 7613
use m3m4contact  m3m4contact_5
timestamp 1652924542
transform -1 0 15785 0 1 5981
box -258 7458 -104 7613
use m3m4contact  m3m4contact_6
timestamp 1652924542
transform -1 0 20049 0 1 6239
box -258 7458 -104 7613
use m3m4contact  m3m4contact_7
timestamp 1652924542
transform -1 0 20049 0 1 5981
box -258 7458 -104 7613
use m3m4contact  m3m4contact_8
timestamp 1652924542
transform 1 0 9789 0 -1 21231
box -258 7458 -104 7613
use m3m4contact  m3m4contact_9
timestamp 1652924542
transform 1 0 9325 0 1 5981
box -258 7458 -104 7613
use m3m4contact  m3m4contact_10
timestamp 1652924542
transform 1 0 13589 0 1 5981
box -258 7458 -104 7613
use m3m4contact  m3m4contact_11
timestamp 1652924542
transform 1 0 14053 0 -1 21231
box -258 7458 -104 7613
use m3m4contact  m3m4contact_12
timestamp 1652924542
transform 1 0 17853 0 1 5981
box -258 7458 -104 7613
use m3m4contact  m3m4contact_13
timestamp 1652924542
transform 1 0 18317 0 -1 21231
box -258 7458 -104 7613
use m3m4contact  m3m4contact_14
timestamp 1652924542
transform 1 0 22117 0 1 5981
box -258 7458 -104 7613
use m3m4contact  m3m4contact_15
timestamp 1652924542
transform 1 0 22581 0 -1 21231
box -258 7458 -104 7613
use m3m4contact  m3m4contact_16
timestamp 1652924542
transform -1 0 8712 0 -1 22211
box -258 7458 -104 7613
use m3m4contact  m3m4contact_17
timestamp 1652924542
transform 1 0 13250 0 -1 22211
box -258 7458 -104 7613
use m3m4contact  m3m4contact_18
timestamp 1652924542
transform -1 0 17240 0 -1 22211
box -258 7458 -104 7613
use m3m4contact  m3m4contact_19
timestamp 1652924542
transform 1 0 21778 0 -1 22211
box -258 7458 -104 7613
use m3m4contact  m3m4contact_20
timestamp 1652924542
transform 1 0 11118 0 -1 22211
box -258 7458 -104 7613
use m3m4contact  m3m4contact_21
timestamp 1652924542
transform 1 0 19646 0 -1 22211
box -258 7458 -104 7613
use m3m4contact  m3m4contact_22
timestamp 1652924542
transform 1 0 11429 0 1 5726
box -258 7458 -104 7613
use m3m4contact  m3m4contact_23
timestamp 1652924542
transform 1 0 19957 0 1 5726
box -258 7458 -104 7613
use m3m4contact  m3m4contact_24
timestamp 1652924542
transform -1 0 11155 0 -1 22917
box -258 7458 -104 7613
use m3m4contact  m3m4contact_25
timestamp 1652924542
transform -1 0 15413 0 -1 22917
box -258 7458 -104 7613
use m3m4contact  m3m4contact_26
timestamp 1652924542
transform 1 0 19957 0 -1 22917
box -258 7458 -104 7613
use m3m4contact  m3m4contact_27
timestamp 1652924542
transform 1 0 15687 0 1 5726
box -258 7458 -104 7613
<< labels >>
flabel metal1 67 695 124 753 0 FreeSans 400 90 0 0 b0
port 1 nsew
flabel metal1 67 2323 124 2381 0 FreeSans 400 0 0 0 b1
port 2 nsew
flabel metal1 67 3951 124 4009 0 FreeSans 400 0 0 0 b2
port 3 nsew
flabel metal1 67 5579 124 5637 0 FreeSans 400 0 0 0 b3
port 4 nsew
flabel metal1 67 7207 124 7265 0 FreeSans 400 0 0 0 b4
port 5 nsew
flabel metal1 67 8835 124 8893 0 FreeSans 400 0 0 0 b5
port 6 nsew
flabel metal1 67 10463 124 10521 0 FreeSans 400 0 0 0 b6
port 7 nsew
flabel metal1 67 12091 124 12149 0 FreeSans 400 0 0 0 b7
port 8 nsew
flabel metal1 63 13539 99 13575 0 FreeSans 320 0 0 0 ena
port 12 nsew
flabel metal3 493 15587 493 15587 0 FreeSans 1600 0 0 0 vss
port 11 nsew
flabel metal4 471 16563 471 16563 0 FreeSans 1600 0 0 0 vdd
port 10 nsew
flabel metal2 234 14816 613 14937 0 FreeSans 1600 0 0 0 dvss
port 14 nsew
flabel metal2 134 14365 427 14487 0 FreeSans 1600 0 0 0 dvdd
port 13 nsew
flabel metal3 7012 121 7012 121 0 FreeSans 480 0 0 0 Vhigh
port 15 nsew
flabel metal3 6588 118 6588 118 0 FreeSans 400 0 0 0 vdd
port 10 nsew
flabel metal3 24656 127 24656 127 0 FreeSans 480 180 0 0 Vlow
port 16 nsew
flabel metal3 24999 118 24999 118 0 FreeSans 400 0 0 0 vss
port 11 nsew
flabel metal4 7332 13732 7332 13732 0 FreeSans 240 0 0 0 b5a
flabel metal4 7332 13477 7332 13477 0 FreeSans 240 0 0 0 b5b
flabel metal3 15545 15638 15545 15638 0 FreeSans 240 90 0 0 out_unbuf
flabel metal2 4570 13896 4570 13896 0 FreeSans 400 90 0 0 b7b
flabel metal2 4722 13892 4722 13892 0 FreeSans 400 90 0 0 b6b
flabel metal2 4875 13893 4875 13893 0 FreeSans 400 90 0 0 b5b
flabel metal2 5024 13895 5024 13895 0 FreeSans 400 90 0 0 b4b
flabel metal2 5179 13898 5179 13898 0 FreeSans 400 90 0 0 b3b
flabel metal2 5328 13897 5328 13897 0 FreeSans 400 90 0 0 b2b
flabel metal2 5483 13885 5483 13885 0 FreeSans 400 90 0 0 b1b
flabel metal2 5634 13897 5634 13897 0 FreeSans 400 90 0 0 b0b
flabel metal2 4647 13897 4647 13897 0 FreeSans 400 90 0 0 b7a
flabel metal2 4799 13896 4799 13896 0 FreeSans 400 90 0 0 b6a
flabel metal2 4952 13892 4952 13892 0 FreeSans 400 90 0 0 b5a
flabel metal2 5103 13894 5103 13894 0 FreeSans 400 90 0 0 b4a
flabel metal2 5256 13896 5256 13896 0 FreeSans 400 90 0 0 b3a
flabel metal2 5406 13897 5406 13897 0 FreeSans 400 90 0 0 b2a
flabel metal2 5560 13885 5560 13885 0 FreeSans 400 90 0 0 b1a
flabel metal2 5711 13892 5711 13892 0 FreeSans 400 90 0 0 b0a
flabel metal3 8596 15634 8596 15634 0 FreeSans 240 180 0 0 b6b
flabel metal3 8715 15638 8715 15638 0 FreeSans 240 180 0 0 b6a
flabel metal3 10851 15638 10851 15638 0 FreeSans 240 180 0 0 b7a
flabel metal3 10726 15638 10726 15638 0 FreeSans 240 180 0 0 b7b
flabel metal3 12861 15634 12861 15634 0 FreeSans 240 180 0 0 b6a
flabel metal3 12975 15634 12975 15634 0 FreeSans 240 180 0 0 b6b
flabel comment 15114 15611 15114 15611 0 FreeSans 240 180 0 0 nca1
flabel comment 14993 15609 14993 15609 0 FreeSans 240 180 0 0 ncb1
flabel metal3 17244 15631 17244 15631 0 FreeSans 240 180 0 0 b6a
flabel metal3 17123 15629 17123 15629 0 FreeSans 240 180 0 0 b6b
flabel metal3 19378 15631 19378 15631 0 FreeSans 240 180 0 0 b7b
flabel metal3 19258 15629 19258 15629 0 FreeSans 240 180 0 0 b7a
flabel metal3 21513 15631 21513 15631 0 FreeSans 240 180 0 0 b6b
flabel metal3 21392 15629 21392 15629 0 FreeSans 240 180 0 0 b6a
flabel comment 23639 15617 23639 15617 0 FreeSans 240 180 0 0 nca2
flabel comment 23518 15615 23518 15615 0 FreeSans 240 180 0 0 ncb2
flabel metal2 16818 21204 17073 21270 0 FreeSans 400 0 0 0 out
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 25939 21270
<< end >>
