magic
tech sky130A
magscale 1 2
timestamp 1652924542
<< metal3 >>
rect -167 7534 -107 7613
rect -169 7528 -105 7534
rect -169 7458 -105 7464
<< via3 >>
rect -169 7464 -105 7528
<< metal4 >>
rect -170 7528 -104 7529
rect -170 7526 -169 7528
rect -258 7466 -169 7526
rect -170 7464 -169 7466
rect -105 7464 -104 7528
rect -170 7463 -104 7464
<< end >>
