magic
tech sky130A
magscale 1 2
timestamp 1652924542
<< xpolycontact >>
rect -35 300 35 732
rect -35 -732 35 -300
<< ppolyres >>
rect -35 -300 35 300
<< viali >>
rect -19 317 19 714
rect -19 -714 19 -317
<< metal1 >>
rect -25 714 25 726
rect -25 317 -19 714
rect 19 317 25 714
rect -25 305 25 317
rect -25 -317 25 -305
rect -25 -714 -19 -317
rect 19 -714 25 -317
rect -25 -726 25 -714
<< res0p35 >>
rect -37 -302 37 302
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 3.0 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 3.854k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
