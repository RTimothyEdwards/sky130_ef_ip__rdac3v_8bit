magic
tech sky130A
magscale 1 2
timestamp 1652995732
<< locali >>
rect 2743 1304 3058 1310
rect 2743 1269 2764 1304
rect 2743 1258 3058 1269
rect 2836 1206 3058 1258
rect 2296 314 2298 367
<< viali >>
rect 2024 1095 2072 1361
rect 3125 1346 4252 1381
rect 2297 1276 2514 1310
rect 2764 1269 4091 1304
rect 3125 1185 4252 1220
rect 481 304 543 438
rect 3151 402 3968 437
rect 2127 314 2296 367
rect 2407 168 2453 345
rect 2845 314 3105 367
rect 3151 241 3968 276
<< metal1 >>
rect 1348 1603 1727 1649
rect -18 1575 1348 1603
rect 1727 1575 4302 1603
rect 3113 1381 4368 1387
rect 2018 1361 2078 1373
rect 2018 1095 2022 1361
rect 2074 1095 2078 1361
rect 3113 1346 3125 1381
rect 4252 1346 4368 1381
rect 3113 1340 4368 1346
rect 2265 1263 2271 1321
rect 2579 1263 2585 1321
rect 2749 1304 4105 1310
rect 2749 1269 2764 1304
rect 4091 1269 4105 1304
rect 2749 1263 4105 1269
rect 3124 1226 3131 1232
rect 3113 1220 3131 1226
rect 3439 1226 3445 1232
rect 4201 1226 4368 1340
rect 3439 1220 4368 1226
rect 3113 1185 3125 1220
rect 4252 1185 4368 1220
rect 3113 1179 3131 1185
rect 3124 1174 3131 1179
rect 3439 1179 4368 1185
rect 3439 1174 3445 1179
rect 2018 1083 2078 1095
rect -18 761 759 863
rect 1138 761 3559 863
rect 3938 761 4302 863
rect 4584 810 4818 874
rect -18 559 220 659
rect 513 559 522 659
rect 4637 651 4695 738
rect 2569 593 4695 651
rect 2569 571 2627 593
rect 1795 513 2627 571
rect 4748 554 4818 810
rect 469 438 555 450
rect 469 401 481 438
rect -17 343 481 401
rect 469 304 481 343
rect 543 401 555 438
rect 1795 401 1853 513
rect 2698 490 4818 554
rect 543 343 1853 401
rect 2016 465 2080 471
rect 543 304 555 343
rect 469 292 555 304
rect 2016 270 2022 465
rect 2074 374 2080 465
rect 2074 367 2308 374
rect 2074 314 2127 367
rect 2296 314 2308 367
rect 2074 308 2308 314
rect 2396 354 2460 357
rect 2074 270 2080 308
rect 2016 264 2080 270
rect 2396 159 2402 354
rect 2454 159 2460 354
rect 2401 156 2459 159
rect -18 21 1348 49
rect 2698 119 2763 490
rect 3139 437 4368 443
rect 3139 402 3151 437
rect 3968 402 4368 437
rect 3139 396 4368 402
rect 2833 370 3117 373
rect 2833 312 2843 370
rect 3107 312 3117 370
rect 2833 308 3117 312
rect 3914 282 4368 396
rect 3139 276 4368 282
rect 3139 241 3151 276
rect 3968 241 4368 276
rect 3139 235 4368 241
rect 1727 21 4302 49
rect 1348 -25 1727 21
<< via1 >>
rect 1348 1501 1727 1603
rect 2022 1095 2024 1361
rect 2024 1095 2072 1361
rect 2072 1095 2074 1361
rect 2271 1310 2579 1321
rect 2271 1276 2297 1310
rect 2297 1276 2514 1310
rect 2514 1276 2579 1310
rect 2271 1263 2579 1276
rect 3131 1220 3439 1232
rect 3131 1185 3439 1220
rect 3131 1174 3439 1185
rect 759 687 1138 937
rect 3559 687 3938 937
rect 220 559 513 659
rect 2022 270 2074 465
rect 2402 345 2454 354
rect 2402 168 2407 345
rect 2407 168 2453 345
rect 2453 168 2454 345
rect 2402 159 2454 168
rect 1348 21 1727 123
rect 2843 367 3107 370
rect 2843 314 2845 367
rect 2845 314 3105 367
rect 3105 314 3107 367
rect 2843 312 3107 314
<< metal2 >>
rect 220 659 513 1669
rect 220 -45 513 559
rect 759 937 1138 1669
rect 759 -45 1138 687
rect 1348 1603 1727 1669
rect 1348 123 1727 1501
rect 2022 1361 2074 1367
rect 2265 1263 2271 1321
rect 2579 1263 2585 1321
rect 2022 465 2074 1095
rect 2022 264 2074 270
rect 2402 354 2454 1263
rect 3124 1174 3131 1232
rect 3439 1174 3445 1232
rect 3138 1062 3229 1174
rect 3007 971 3229 1062
rect 3007 370 3098 971
rect 3559 937 3938 1669
rect 2837 312 2843 370
rect 3107 312 3113 370
rect 2402 153 2454 159
rect 1348 -50 1727 21
rect 3559 -45 3938 687
use sky130_fd_pr__diode_pw2nd_05v5_4AXGXB  sky130_fd_pr__diode_pw2nd_05v5_4AXGXB_0 paramcells
timestamp 1652928066
transform 1 0 4664 0 1 721
box -183 -183 183 183
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1650294714
transform 1 0 4206 0 1 -2
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1650294714
transform 1 0 4014 0 1 -2
box -66 -43 258 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1650294714
transform 1 0 2094 0 1 -2
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1650294714
transform 1 0 2094 0 -1 1626
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_8  sky130_fd_sc_hvl__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1650294714
transform 1 0 2862 0 -1 1626
box -66 -43 1506 897
use sky130_fd_sc_hvl__inv_8  sky130_fd_sc_hvl__inv_8_1
timestamp 1650294714
transform 1 0 2574 0 1 -2
box -66 -43 1506 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1650294714
transform 1 0 -18 0 1 -2
box -66 -43 2178 1671
<< labels >>
flabel metal1 194 372 194 372 0 FreeSans 480 0 0 0 bit_in
flabel metal1 174 609 174 609 0 FreeSans 480 0 0 0 dvdd
flabel metal2 938 1039 938 1039 0 FreeSans 480 0 0 0 avdd
flabel metal2 1508 1392 1508 1392 0 FreeSans 480 0 0 0 agnd
flabel metal2 3738 1039 3738 1039 0 FreeSans 480 0 0 0 avdd
flabel metal1 4287 331 4287 331 0 FreeSans 480 0 0 0 bit_out
flabel metal1 4276 1286 4276 1286 0 FreeSans 480 0 0 0 bitb_out
<< end >>
