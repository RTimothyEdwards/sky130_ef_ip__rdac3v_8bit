magic
tech sky130A
magscale 1 2
timestamp 1652924542
<< nwell >>
rect 316 892 942 1410
rect 318 -275 942 228
<< mvpsubdiff >>
rect 573 590 687 595
rect 573 530 599 590
rect 663 530 687 590
rect 573 525 687 530
<< mvnsubdiff >>
rect 496 1298 520 1344
rect 743 1298 767 1344
rect 496 -209 520 -163
rect 743 -209 767 -163
<< mvpsubdiffcont >>
rect 599 530 663 590
<< mvnsubdiffcont >>
rect 520 1298 743 1344
rect 520 -209 743 -163
<< locali >>
rect 496 1298 520 1344
rect 743 1298 767 1344
rect 599 590 664 606
rect 599 514 664 530
rect 496 -209 520 -163
rect 743 -209 767 -163
<< viali >>
rect 613 1298 652 1301
rect 613 1222 652 1298
rect 599 530 663 590
rect 663 530 664 590
rect 613 -163 652 -85
rect 613 -166 652 -163
<< metal1 >>
rect 600 1307 665 1322
rect 290 1199 446 1245
rect 600 1215 606 1307
rect 659 1215 665 1307
rect 992 1284 1105 1339
rect 600 1209 665 1215
rect 814 1199 960 1245
rect 290 1176 342 1199
rect 290 1114 342 1124
rect 908 1046 960 1199
rect 908 984 960 994
rect 390 911 436 958
rect 548 911 594 958
rect 666 911 712 958
rect 387 905 439 911
rect 387 847 439 853
rect 545 905 597 911
rect 545 847 597 853
rect 663 905 715 911
rect 663 847 715 853
rect 824 896 870 958
rect 992 896 1026 1284
rect 824 862 1026 896
rect 290 807 342 813
rect 390 799 436 847
rect 548 799 594 847
rect 666 799 712 847
rect 824 799 870 862
rect 290 637 342 755
rect 918 789 970 795
rect 918 637 970 737
rect 290 591 446 637
rect 604 609 659 615
rect 593 590 604 602
rect 659 590 671 602
rect 814 591 970 637
rect 593 530 599 590
rect 664 530 671 590
rect 290 483 446 529
rect 593 518 604 530
rect 659 518 671 530
rect 604 506 659 512
rect 814 483 970 529
rect 290 402 342 483
rect 290 344 342 350
rect 918 383 970 483
rect 918 325 970 331
rect 390 258 436 321
rect 548 276 594 321
rect 666 276 712 321
rect 824 276 870 321
rect 234 224 436 258
rect 234 -168 268 224
rect 390 162 436 224
rect 545 270 597 276
rect 545 212 597 218
rect 663 270 715 276
rect 663 212 715 218
rect 821 270 873 276
rect 821 212 873 218
rect 548 162 594 212
rect 666 162 712 212
rect 824 162 870 212
rect 300 142 352 148
rect 300 -79 352 90
rect 918 16 970 22
rect 600 -78 665 -72
rect 300 -125 446 -79
rect 155 -223 268 -168
rect 600 -172 606 -78
rect 659 -172 665 -78
rect 918 -79 970 -36
rect 814 -125 970 -79
rect 600 -185 665 -172
<< via1 >>
rect 606 1301 659 1307
rect 606 1222 613 1301
rect 613 1222 652 1301
rect 652 1222 659 1301
rect 606 1215 659 1222
rect 290 1124 342 1176
rect 908 994 960 1046
rect 387 853 439 905
rect 545 853 597 905
rect 663 853 715 905
rect 290 755 342 807
rect 918 737 970 789
rect 604 590 659 609
rect 604 530 659 590
rect 604 512 659 530
rect 290 350 342 402
rect 918 331 970 383
rect 545 218 597 270
rect 663 218 715 270
rect 821 218 873 270
rect 300 90 352 142
rect 918 -36 970 16
rect 606 -85 659 -78
rect 606 -166 613 -85
rect 613 -166 652 -85
rect 652 -166 659 -85
rect 606 -172 659 -166
<< metal2 >>
rect 99 1307 1166 1347
rect 99 1215 606 1307
rect 659 1215 1166 1307
rect 99 1210 1166 1215
rect 144 1122 153 1178
rect 209 1176 218 1178
rect 209 1124 290 1176
rect 342 1124 348 1176
rect 209 1122 218 1124
rect 1043 1046 1052 1048
rect 902 994 908 1046
rect 960 994 1052 1046
rect 1043 992 1052 994
rect 1108 992 1117 1048
rect 376 905 450 907
rect 376 853 387 905
rect 439 853 450 905
rect 376 851 450 853
rect 529 905 608 907
rect 529 853 545 905
rect 597 853 608 905
rect 529 851 608 853
rect 652 905 729 907
rect 652 853 663 905
rect 715 853 729 905
rect 652 851 729 853
rect 143 753 152 809
rect 208 807 217 809
rect 208 755 290 807
rect 342 755 348 807
rect 1043 789 1052 791
rect 208 753 217 755
rect 912 737 918 789
rect 970 737 1052 789
rect 1043 735 1052 737
rect 1108 735 1117 791
rect 99 609 1166 678
rect 99 512 604 609
rect 659 512 1166 609
rect 99 453 1166 512
rect 143 348 152 404
rect 208 402 217 404
rect 208 350 290 402
rect 342 350 348 402
rect 1043 383 1052 385
rect 208 348 217 350
rect 912 331 918 383
rect 970 331 1052 383
rect 1043 329 1052 331
rect 1108 329 1117 385
rect 529 270 608 272
rect 529 218 545 270
rect 597 218 608 270
rect 529 216 608 218
rect 652 270 731 273
rect 652 218 663 270
rect 715 218 731 270
rect 652 217 731 218
rect 810 270 883 272
rect 810 218 821 270
rect 873 218 883 270
rect 810 216 883 218
rect 143 88 152 144
rect 208 142 217 144
rect 208 90 300 142
rect 352 90 358 142
rect 208 88 217 90
rect 1044 16 1053 18
rect 912 -36 918 16
rect 970 -36 1053 16
rect 1044 -38 1053 -36
rect 1109 -38 1118 18
rect 99 -78 1166 -72
rect 99 -172 606 -78
rect 659 -172 1166 -78
rect 99 -210 1166 -172
<< via2 >>
rect 153 1122 209 1178
rect 1052 992 1108 1048
rect 152 753 208 809
rect 1052 735 1108 791
rect 152 348 208 404
rect 1052 329 1108 385
rect 152 88 208 144
rect 1053 -38 1109 18
<< metal3 >>
rect 148 1178 214 1188
rect 148 1122 153 1178
rect 209 1122 214 1178
rect 148 1121 214 1122
rect 148 1057 149 1121
rect 213 1057 214 1121
rect 148 1038 214 1057
rect 1047 1048 1113 1058
rect 1047 992 1052 1048
rect 1108 992 1113 1048
rect 1047 928 1048 992
rect 1112 928 1113 992
rect 1047 908 1113 928
rect 147 863 213 882
rect 147 799 148 863
rect 212 799 213 863
rect 147 753 152 799
rect 208 753 213 799
rect 147 731 213 753
rect 1047 791 1113 801
rect 1047 735 1052 791
rect 1108 735 1113 791
rect 1047 734 1113 735
rect 1047 670 1048 734
rect 1112 670 1113 734
rect 1047 651 1113 670
rect 147 467 213 488
rect 147 403 148 467
rect 212 403 213 467
rect 147 348 152 403
rect 208 348 213 403
rect 147 338 213 348
rect 1047 385 1113 393
rect 1047 338 1052 385
rect 1108 338 1113 385
rect 1047 274 1048 338
rect 1112 274 1113 338
rect 1047 241 1113 274
rect 147 208 213 228
rect 147 144 148 208
rect 212 144 213 208
rect 147 88 152 144
rect 208 88 213 144
rect 147 78 213 88
rect 1048 82 1114 102
rect 1048 18 1049 82
rect 1113 18 1114 82
rect 1048 -38 1053 18
rect 1109 -38 1114 18
rect 1048 -48 1114 -38
<< via3 >>
rect 149 1057 213 1121
rect 1048 928 1112 992
rect 148 809 212 863
rect 148 799 152 809
rect 152 799 208 809
rect 208 799 212 809
rect 1048 670 1112 734
rect 148 404 212 467
rect 148 403 152 404
rect 152 403 208 404
rect 208 403 212 404
rect 1048 329 1052 338
rect 1052 329 1108 338
rect 1108 329 1112 338
rect 1048 274 1112 329
rect 148 144 212 208
rect 1049 18 1113 82
<< metal4 >>
rect 148 1121 214 1122
rect 148 1119 149 1121
rect 99 1059 149 1119
rect 148 1057 149 1059
rect 213 1119 214 1121
rect 213 1059 1166 1119
rect 213 1057 214 1059
rect 148 1056 214 1057
rect 1047 992 1113 993
rect 1047 990 1048 992
rect 99 930 1048 990
rect 1047 928 1048 930
rect 1112 990 1113 992
rect 1112 930 1166 990
rect 1112 928 1113 930
rect 1047 927 1113 928
rect 147 863 213 864
rect 147 861 148 863
rect 99 801 148 861
rect 147 799 148 801
rect 212 861 213 863
rect 212 801 1166 861
rect 212 799 213 801
rect 147 798 213 799
rect 1047 734 1113 735
rect 1047 732 1048 734
rect 99 672 1048 732
rect 1047 670 1048 672
rect 1112 732 1113 734
rect 1112 672 1166 732
rect 1112 670 1113 672
rect 1047 669 1113 670
rect 147 467 213 468
rect 147 465 148 467
rect 99 405 148 465
rect 147 403 148 405
rect 212 465 213 467
rect 212 405 1166 465
rect 212 403 213 405
rect 147 402 213 403
rect 1047 338 1113 339
rect 1047 336 1048 338
rect 99 276 1048 336
rect 1047 274 1048 276
rect 1112 336 1113 338
rect 1112 276 1166 336
rect 1112 274 1113 276
rect 1047 273 1113 274
rect 147 208 213 209
rect 147 207 148 208
rect 99 147 148 207
rect 147 144 148 147
rect 212 207 213 208
rect 212 147 1166 207
rect 212 144 213 147
rect 147 143 213 144
rect 1048 82 1114 83
rect 1048 78 1049 82
rect 99 18 1049 78
rect 1113 78 1114 82
rect 1113 18 1166 78
rect 1048 17 1114 18
use sky130_fd_pr__nfet_g5v0d10v5_NHLDUY  sky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 paramcells
timestamp 1652924542
transform 1 0 492 0 1 703
box -108 -122 108 122
use sky130_fd_pr__nfet_g5v0d10v5_NHLDUY  sky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1
timestamp 1652924542
transform 1 0 768 0 1 703
box -108 -122 108 122
use sky130_fd_pr__nfet_g5v0d10v5_NHLDUY  sky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2
timestamp 1652924542
transform 1 0 492 0 -1 417
box -108 -122 108 122
use sky130_fd_pr__nfet_g5v0d10v5_NHLDUY  sky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3
timestamp 1652924542
transform 1 0 768 0 -1 417
box -108 -122 108 122
use sky130_fd_pr__pfet_g5v0d10v5_9992MR  sky130_fd_pr__pfet_g5v0d10v5_9992MR_0 paramcells
timestamp 1652924542
transform 1 0 492 0 1 1094
box -174 -202 174 164
use sky130_fd_pr__pfet_g5v0d10v5_9992MR  sky130_fd_pr__pfet_g5v0d10v5_9992MR_1
timestamp 1652924542
transform 1 0 768 0 1 1094
box -174 -202 174 164
use sky130_fd_pr__pfet_g5v0d10v5_9992MR  sky130_fd_pr__pfet_g5v0d10v5_9992MR_2
timestamp 1652924542
transform 1 0 768 0 -1 26
box -174 -202 174 164
use sky130_fd_pr__pfet_g5v0d10v5_9992MR  sky130_fd_pr__pfet_g5v0d10v5_9992MR_3
timestamp 1652924542
transform 1 0 492 0 -1 26
box -174 -202 174 164
use sky130_fd_pr__res_high_po_0p35_AW5QUD  sky130_fd_pr__res_high_po_0p35_AW5QUD_0 paramcells
timestamp 1652924542
transform 1 0 180 0 1 558
box -37 -732 37 732
use sky130_fd_pr__res_high_po_0p35_AW5QUD  sky130_fd_pr__res_high_po_0p35_AW5QUD_1
timestamp 1652924542
transform 1 0 1080 0 1 558
box -37 -732 37 732
<< end >>
